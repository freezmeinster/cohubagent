module command

import cli { Command, Flag }

pub fn list_func(cmd Command) {
    println("cuk")
}
